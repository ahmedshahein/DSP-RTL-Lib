/home/shahein/ENGINEERING/CODES/verilog/ppd/dsp_filt_mac/sim/testcases/stimuli/defines_9.sv