/home/shahein/ENGINEERING/CODES/verilog/dsp_rtl_lib/filt_ppi/sim/testcases/stimuli/defines_4.sv