`define P_INP_W 	8
`define P_OUP_W 	16
`define P_FF_COEF_L 	3
`define P_FF_COEFF_W 	8
`define P_FB_COEFF_L 	3
`define P_FB_COEFF_W 	8
`define P_TOPOLOGY 	0

`define TESTCASE	1

`define NULL 	0