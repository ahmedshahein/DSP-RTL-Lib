/home/shahein/ENGINEERING/CODES/verilog/ppd/dsp_filt_ppi/sim/testcases/stimuli/defines_5.sv