`define P_INP_DATA_W 	2
`define P_COEFF_L 	32
`define P_COEFF_W 	16
`define P_SYMM 		0
`define P_OUP_DATA_W 	50

`define TESTCASE	3

`define DIV2(N) ((N/2)+(N%2))

`define NULL 	0