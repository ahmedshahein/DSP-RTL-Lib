`define DIV(N, D) (N%D==0) ? (N/D) : (N/D+1)

`define P_INP_DATA_W 	6
`define P_DECIMATION 	31
`define P_COEFF_L 	53
`define P_COEFF_W 	16
`define P_TF_DF 	1
`define P_COMM_R_OUP 	1
`define P_COMM_CCW_CW 	1
`define P_MUL_CCW_CW 	0
`define P_COMM_PHA 	0
`define P_OUP_W     	28

`define TESTCASE	8

`define NULL 	0