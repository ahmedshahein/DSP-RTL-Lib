`define P_ROM_WIDTH 		16
`define P_ROM_DEPTH 		13
`define P_PHASEACCU_WIDTH 	32

`define TESTCASE		4

`define NULL 	0