`define P_INTERPOLATION 13
`define P_ORDER 	5
`define P_DIFF_DELAY 	1
`define P_PHASE 	7
`define P_INP_DATA_W 	8
`define P_OUP_DATA_W 	28

`define TESTCASE	8

`define NULL 	0