`define P_DECIMATION 	16
`define P_ORDER 	8
`define P_DIFF_DELAY 	1
`define P_PHASE 	3
`define P_INP_DATA_W 	2
`define P_OUP_DATA_W 	34

`define TESTCASE	3

`define NULL 	0