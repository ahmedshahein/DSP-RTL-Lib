`define P_INP_DATA_W 	8
`define P_COEFF_L 	33
`define P_COEFF_W 	12
`define P_TF_DF 	1
`define P_SYMM 		1
`define P_OUP_DATA_W 	53

`define TESTCASE	3

`define NULL 	0