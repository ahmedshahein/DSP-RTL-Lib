/home/shahein/ENGINEERING/CODES/verilog/ppd/dsp_filt_ppd/sim/testcases/stimuli/defines_5.sv