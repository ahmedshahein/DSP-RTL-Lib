`define P_DECIMATION 	32
`define P_ORDER 	5
`define P_DIFF_DELAY 	1
`define P_PHASE 	0
`define P_INP_DATA_W 	8
`define P_OUP_DATA_W 	33

`define TESTCASE	1

`define NULL 	0