/home/shahein/ENGINEERING/CODES/verilog/dsp_rtl_lib/filt_cici/sim/testcases/stimuli/defines_7.sv