/home/shahein/ENGINEERING/CODES/verilog/ppd/dsp_nco/sim/testcases/stimuli/defines_4.sv