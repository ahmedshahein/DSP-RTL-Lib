/home/shahein/ENGINEERING/CODES/verilog/dsp_rtl_lib/filt_cic/sim/testcases/stimuli/defines_1.sv