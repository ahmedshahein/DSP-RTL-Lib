`define P_INP_DATA_W 	7
`define P_COEFF_L 	64
`define P_COEFF_W 	13
`define P_TF_DF 	0
`define P_SYMM 		1
`define P_OUP_DATA_W 	26

`define TESTCASE	9

`define NULL 	0