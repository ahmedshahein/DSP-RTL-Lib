/home/shahein/ENGINEERING/CODES/verilog/dsp_rtl_lib/filt_mac/sim/testcases/stimuli/defines_5.sv