/home/shahein/ENGINEERING/CODES/verilog/dsp_rtl_lib/filt_ppd/sim/testcases/stimuli/defines_9.sv