/home/shahein/ENGINEERING/CODES/verilog/dsp_rtl_lib/sgen_nco/sim/testcases/stimuli/defines_1.sv