/home/shahein/ENGINEERING/CODES/verilog/ppd/dsp_filt_fir/sim/testcases/stimuli/defines_1.sv